netcdf PCASP1_cal_template {

// This cdl file contains the attributes, dimensions, and variables that are
// applied to all calibration netCDF files for a particular instrument.
//
// Instrument: PCASP-1
//
// Structure of the cal-nc file is as follows ;
// Global attributes
//  Group: bin_cal
//      Contains scattering cross-section calibration info for size bins.
//    Group: Secondary material sub-group
//      This sub-group of bin_cal/ contains diameter-related variables for
//      another material. Dimensions are inherited from bin_cal. Material
//      information is included in group and variable attributes.
//    Group: Another material sub-group
//      Any number of material sub-groups can be included for different
//      particle types/materials.
//
// author = G. Nott
// email = graeme.nott@faam.ac.uk
// creation = Jan 2021

// global attributes:

    // Universal global file attributes. Do not modify.
    :Conventions = "CF-1.7" ;
    :_Format = "netCDF-4" ;
    :institution = "FAAM. Facility for Airborne Atmospheric Measurements" ;
    :address = "Building 146, Cranfield University, Cranfield MK43 0AL UK" ;
    :software_repository = "https://github.com/FAAM-146/cal-nc" ;

    // Instrument global file attributes.
    :title = "FAAM calibration data for the PCASP-1" ;
    :source = "Laboratory-based calibration" ;
    :instr = "PCASP-1" ;
    :instr_long_name = "Passive Cavity Spectrometer Probe. SPP200 electronics package" ;
    :instr_serialnumber = "17884-0190-04" ;
    :references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;

// The following global attributes shall be modified by cal_ncgen.py if used
    :username = ;
    :history = ;


group: bin_cal {
    // Group containing calibration of size bins of the PCASP

    :title = "Size bin calibration of PCASP" ;
    :comment = "Group containing calibration of size bins of the PCASP. Photodetector voltage pulse-heights are calibrated to the calculated scattering cross-section of known PSL and DEHS monodisperse distributions." ;
    :references = "P.D. Rosenberg, A.R. Dean, P.I. Williams, J.R. Dorsey, A. Minikin, M.A. Pickering and A. Petzold, Particle sizing calibration with refractive index correction for light scattering optical particle counters and impacts upon PCASP and CDP data collected during the Fennec campaign, Atmos. Meas. Tech., 5, 1147-1163, doi:10.5194/amt-5-1147-2012, 2012." ;
    :applied = "False" ;

    // Define dimensions for group.
    dimensions:
        time = UNLIMITED ;
        bin = 30 ;
        bin_bounds = 2 ;

    // Define group coordinate variable
    variables:
        float time(time) ;
            // The units of time may be one of days ('d'), hours ('hr', 'h'),
            // minutes ('min'), or seconds ('sec', 's'). The most appropriate
            // unit given the frequency of calibration should be used.
            time:standard_name = "time" ;
            time:long_name = "time of calibration" ;
            time:timezone = "UTC" ;
            time:units = "seconds since 1970-01-01 00:00:00" ;
            time:strftime_format = "seconds since %Y-%m-%d %H:%M:%S%Z" ;

        int bin(bin) ;
            bin:long_name = "bin number" ;
            bin:comment = "The PCASP has 30 bins however the first has a somewhat undefined lower boundary and should therefore usually be discarded." ;

    // Define group variables
        string applies_to(time) ;
            applies_to:long_name = "Calibration applies to this data" ;
            applies_to:comment = "String of applicable flight numbers or other unique identifier for each calibration time/date" ;

        string descr(time) ;
            descr:long_name = "Description of calibration" ;
            descr:comment = "Any descriptive string used as an addition identifier of this calibration" ;

        string traceability(time) ;
            traceability:long_name = "Traceability of calibration" ;
            traceability:comment = "Link to file/s showing traceability of calibration materials and instruments or unique lot numbers for each calibration PSL." ;

        string calibration_file(time) ;
            calibration_file:long_name = "File from which this calibration data has been read" ;

        string source_file(time) ;
            source_file:long_name = "Source file used in calibration processing" ;

        int cal_flag(time) ;
            cal_flag:long_name = "Flag denoting quality of calibration" ;
            cal_flag:valid_range = 0, 3 ;
            cal_flag:flag_values = 0, 1, 2, 3 ;
            cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
            cal_flag:_FillValue = 3 ;

        int ADC_thres(time,bin,bin_bounds) ;
            ADC_thres:long_name = "Lower and upper ADC thresholds for each bin" ;
            ADC_thres:comment = "Coverage of each bin in terms of the digitized peak photovoltage. This variable has been included primarily for error checking as the same values should be in the standard data files." ;
            ADC_thres:valid_range = 0, 12288 ;
            ADC_thres:_FillValue = NaN ;

        float x-section(time,bin,bin_bounds) ;
            x-section:long_name = "Lower and upper scattering cross-section boundaries for each bin" ;
            x-section:comment = "Lower boundary of first bin is undefined." ;
            x-section:units = "um**2" ;
            x-section:ancillary_variables = "x-section_err" ;
            x-section:_FillValue = NaN ;

        float x-section_err(time,bin,bin_bounds) ;
            x-section_err:long_name = "Uncertainty of scattering cross-section boundaries for each bin" ;
            x-section_err:comment = "Uncertainties are derived from the uncertainty in the calculated scattering cross-section and the width of the modal bin for each calibration particle. These are discussed in sections 2.1 and 2.23 in Rosenberg et al. (full citation given in references attribute of this group)." ;
            x-section_err:_FillValue = NaN ;

        float x-section_width(time,bin) ;
            x-section_width:long_name = "Width of each bin in terms of scattering cross-section" ;
            x-section:units = "um**2" ;
            x-section:ancillary_variables = "x-section_width_err" ;
            x-section:_FillValue = NaN ;

        float x-section_width_err(time,bin) ;
            x-section_width_err:long_name = "Uncertainty of scattering cross-section width for each bin" ;
            x-section_width_err:comment = "Uncertainties are derived from the uncertainty in the calculated scattering cross-section and the width of the modal bin for each calibration particle. These are discussed in sections 2.1 and 2.23 in Rosenberg et al. (full citation given in references attribute of this group)." ;
            x-section_width_err:_FillValue = NaN ;


    data:
        // Data is comma-delineated with no additional deliniation between
        // dimensions. Thus the data is presented flattened with the overall
        // length being d1*d2*..dn. As specified in the variable definition,
        // the dimensions are cycled over in reverse order so for multi-
        // dimensional arrays, the last dimension varies fastest. Thus,
        // row-order rather than column order is used for matrices. If
        // var = np.array([[11,12,13],[21,22,23]]) then var.flatten() or
        // np.ravel(var) will write the array in the correct way.
        // Missing data can be written as '_'

        bin = 1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30 ;


    group: mineral_dust {
        // Group containing calibration of size bins of the PCASP for mineral dust

        // MOVE THIS TO SEPARATE CDL FILE IN DATA DIR
        // HMM, CAN THIS BE DONE WITH PARENT COORDS?


        :title = "Size bin diameter calibrations of PCASP for mineral dust" ;
        :comment = "The real part of the refractive index was taken as 1.53 which is a common value and is in the OPAC database. It is quite a bit smaller than the 1.547 that was reported by Weinzierl et al. [2011] but has been shown to have a relatively weak effect on the instrument response. The values of the imaginary part were based on references in  Ryder et al. [2019] along with the frequency distribution of k(550nm) presented in fig 9 of Ryder et al. [2013]. So the minimum value was extended from 0.0015i to 0.001i. Calculating the bin boundaries with these multiple Mie curves was done with Gaussian centre-weighted averaging with 0.001i and 0.0024i being +/-2 sigma extreme values." ;
        :references = "Weinzierl et al., Tellus 63B, 589-618, 2011., Ryder et al., ACP 19, 5353-15376, 2019, Ryder et al., ACP 13, 303-325, 2013." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float dia_centre(time,bin) ;
                dia_centre:long_name = "Centre diameter of each bin for given particle material - mineral dust" ;
                dia_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. (full citation given in references attribute of this group)." ;
                dia_centre:refractive_index = "1.53 + (0.001i--0.0024i)" ;
                dia_centre:shape = "spherical" ;
                dia_centre:units = "um" ;
                dia_centre:ancillary_variables = "dia_centre_err dia_width" ;
                dia_centre:_FillValue = NaN ;

            float dia_centre_err(time,bin) ;
                dia_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                dia_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                dia_centre_err:units = "um" ;
                dia_centre_err:_FillValue = NaN ;

            float dia_width(time,bin) ;
                dia_width:long_name = "Width in terms of diameter of each bin for given particle material - mineral dust" ;
                dia_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                dia_width:refractive_index = "1.53 + (0.001i--0.0024i)" ;
                dia_width:shape = "spherical" ;
                dia_width:units = "um" ;
                dia_width:ancillary_variables = "dia_width_err" ;
                dia_width:_FillValue = NaN ;

            float dia_width_err(time,bin) ;
                dia_width_err:long_name = "Uncertainty of bin diameter width" ;
                dia_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                dia_width_err:units = "um" ;
                dia_width_err:_FillValue = NaN ;

        } // End group bin_cal/mineral_dust

    } // End group bin_cal


group: flow_cal {
    // Group containing calibration of flow rates of the PCASP
    //
    :title = "Flow calibration of PCASP" ;
    :comment = "Group containing sample flow calibration information. Sample flow output and/or input is measured by a calibrated meter" ;
    :references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
    :applied = "True" ;

    // The units of time may be one of days ('d'), hours ('hr', 'h'),
    // minutes ('min'), or seconds ('sec', 's') and the most appropriate unit
    // for the frequency of calibration should be used.
    dimensions:
        time = UNLIMITED ;
        max_flows = 32 ;    // Maximum number of different flows in a calibration

    // Define group coordinate variable
    variables:
        float time(time) ;
            // The units of time may be one of days ('d'), hours ('hr', 'h'),
            // minutes ('min'), or seconds ('sec', 's') and the most appropriate
            // unit for the frequency of calibration should be used.
            time:standard_name = "time" ;
            time:long_name = "time of calibration" ;
            time:timezone = "UTC" ;
            time:units = "seconds since 1970-01-01 00:00:00" ;
            time:strftime_format = "seconds since %Y-%m-%d %H:%M:%S%Z" ;

    // Define group variables
        string applies_to(time) ;
            applies_to:long_name = "Calibration applies to this data" ;
            applies_to:comments = "String of applicable flight numbers or other unique identifier for calibration." ;

        string descr(time) ;
            descr:long_name = "Description of calibration" ;
            descr:comment = "Any descriptive string used as an addition identifier of this calibration." ;

        string traceability(time) ;
            traceability:long_name = "Traceability of calibration" ;
            traceability:comment = "Links to calibration certificates or other identifiers showing traceability of calibration instruments." ;

        int cal_flag(time) ;
            cal_flag:long_name = "Flag denoting quality of calibration" ;
            cal_flag:valid_range = 0, 3 ;
            cal_flag:flag_values = 0, 1, 2, 3 ;
            cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
            cal_flag:_FillValue = 3 ;

        float flows_reported(time,max_flows) ;
            flows_reported:long_name = "Sample flow rate reported by PCASP for each value in flows_actual" ;
            flows_reported:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the length of flows_reported for each time is the same as flows_actual for that time." ;
            flows_reported:units = "cc/s" ;
//            flows_reported:valid_min = -0.01 ;
            flows_reported:_FillValue = NaN ;

        float flows_actual(time,max_flows) ;
            flows_actual:long_name = "Verified sample flow rate for each value in flows_reported" ;
            flows_actual:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_actual for each time is the same as flows_reported for that time." ;
            flows_actual:units = "cc/s" ;
//            flows_actual:valid_min = -0.01 ;
            flows_actual:_FillValue = NaN ;

        string flow_fit(time) ;
            flow_fit:long_name = "Calibration equation of sample flow" ;
            flow_fit:comment = "String of equation used to convert reported sample flow to calibrated sample flow rate. This will involve a fit to the data given for the same time stamp in the flows variable. A string is used for flexibility but may be changed to polynomial values in the future if appropriate." ;
        flow_fit:_FillValue = "" ;


    data:
        // Data is comma-delineated with no additional deliniation between
        // dimensions. Thus the data is presented flattened with the overall
        // length being d1*d2*..dn. As specified in the variable definition,
        // the dimensions are cycled over in reverse order so for multi-
        // dimensional arrays, the last dimension varies fastest. Thus,
        // row-order rather than column order is used for matrices.. If
        // var = np.array([[11,12,13],[21,22,23]]) then var.flatten() or
        // np.ravel(var) will write the array in the correct way.

    } // End group flow_cal

} // EOF