netcdf \20191107_P2_cal {

// global attributes:
		:Conventions = "CF-1.6" ;
		:NCO = "4.1.3" ;
		:institution = "FAAM. Facility for Airborne Atmospheric Measurements" ;
		:address = "Building 146, Cranfield University, Cranfield MK43 0AL UK" ;
		:title = "FAAM calibration data for the PCASP-2" ;
		:source = "Laboratory-based calibration" ;
		:instr = "PCASP-2" ;
		:instr_long_name = "Passive Cavity Spectrometer Probe. SPP200 electronics package" ;
		:instr_serialnumber = "PMI-1022-1202-31" ;
		:references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
		:username = "Graeme Nott <graeme.nott@faam.ac.uk>" ;
		:history = "20191129T0957 Initial creation" ;
		:software_version = "0.2" ;

group: bin_cal {
  dimensions:
  	time = UNLIMITED ; // (2 currently)
  	bin = 30 ;
  	bin_bounds = 2 ;
  variables:
  	float time(time) ;
  		time:standard_name = "time" ;
  		time:long_name = "time of calibration" ;
  		time:timezone = "UTC" ;
  		time:units = "days since 1970-01-01 00:00:00" ;
  		time:strftime_format = "days since %Y-%m-%d %Z" ;
  	int bin(bin) ;
  		bin:long_name = "bin number" ;
  		bin:comment = "The PCASP has 30 bins however the first has a somewhat undefined lower boundary and should therefore usually be discarded." ;
  	string applies_to(time) ;
  		applies_to:long_name = "Each calibration applies to these measurements" ;
  		applies_to:comment = "String of applicable flight numbers for calibration" ;
  	string descr(time) ;
  		descr:long_name = "Description of calibration" ;
  		descr:comment = "Campaign name/s for which these calibrations apply" ;
  	string traceability(time) ;
  		traceability:long_name = "Traceability trail for each calibration" ;
  		traceability:comment = "Unique lot numbers for each calibration PSL. These can be traced to the original NIST-traceable certificates." ;
  	int cal_flag(time) ;
  		cal_flag:long_name = "Flag denoting quality of calibration" ;
  		cal_flag:valid_range = 0, 3 ;
  		cal_flag:flag_values = 0, 1, 2, 3 ;
  		cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
  		cal_flag:_FillValue = 3 ;
  	int ADC_thres(time, bin, bin_bounds) ;
  		ADC_thres:long_name = "Lower and upper ADC thresholds for each bin" ;
  		ADC_thres:comment = "Coverage of each bin in terms of the digitized peak photovoltage. This variable has been included primarily for error checking as the same values should be in the standard data files." ;
  		ADC_thres:valid_range = 0, 12289 ;
  		ADC_thres:_FillValue = -2147483648 ;
  	float x-section(time, bin, bin_bounds) ;
  		x-section:long_name = "Scattering cross-section boundaries for each bin" ;
  		x-section:comment = "Lower boundary of first bin is undefined." ;
  		x-section:units = "m**2" ;
  		x-section:ancillary_variables = "x-section_width_err" ;
  		x-section:_FillValue = -9999.f ;
  	float x-section_err(time, bin, bin_bounds) ;
  		x-section_err:long_name = "Uncertainty of scattering cross section boundaries for each bin" ;
  		x-section_err:comment = "Straight-line fits for scattering cross-section versus ADC voltage are calculated along with sensitivities to the uncertainty in these data. See section 2.2.3 of Rosenberg et al. (2012) for details." ;
  		x-section_err:_FillValue = -9999.f ;
  	float x-section_width(time, bin) ;
  		x-section_width:long_name = "Width of each bin in terms of scattering cross section" ;
  	float x-section_width_err(time, bin) ;
  		x-section_width_err:long_name = "Uncertainty of scattering cross section boundaries for each bin" ;
  		x-section_width_err:comment = "" ;
  		x-section_width_err:flag_values = 0, 1 ;
  		x-section_width_err:flag_meanings = "Independent_uncertainties \n                                                 Dependent_uncertainties" ;
  		x-section_width_err:_FillValue = -9999.f ;
  	float dia_centre(time, bin) ;
  		dia_centre:long_name = "Centre diameter associated with each bin number for given particle material properties" ;
  		dia_centre:comment = "This is the weighted average of each of the regions of the scattering curve which include the range of scattering cross-sections in each bin with the uncertainty of these boundaries included. This is discussed in sections 4.1 and 4.2 of Rosenberg et al. (2012)." ;
  		dia_centre:refractive_index = "1.59+0i" ;
  		dia_centre:shape = "spherical" ;
  		dia_centre:units = "um" ;
  		dia_centre:ancillary_variables = "dia_centre_err dia_width" ;
  		dia_centre:_FillValue = -9999.f ;
  	float dia_centre_err(time, bin) ;
  		dia_centre_err:long_name = "Uncertainty of bin centre diameter" ;
  		dia_centre_err:comment = "See sections 4.1 and 4.2 of Rosenberg et al. (2012). for details." ;
  		dia_centre_err:units = "um" ;
  		dia_centre_err:_FillValue = -9999.f ;
  	float dia_width(time, bin) ;
  		dia_width:long_name = "Diameter width associated with each bin number for given particle material properties" ;
  		dia_width:comment = "This is the sum of all regions of the scattering curve which include the range of scattering cross-sections in each bin with the uncertainty of these boundaries included. This is discussed in sections 4.1 and 4.2 of Rosenberg et al. (2012)." ;
  		dia_width:refractive_index = "1.59+0i" ;
  		dia_width:shape = "spherical" ;
  		dia_width:units = "um" ;
  		dia_width:ancillary_variables = "dia_width_err" ;
  		dia_width:_FillValue = -9999.f ;
  	float dia_width_err(time, bin) ;
  		dia_width_err:long_name = "Uncertainty of bin width" ;
  		dia_width_err:comment = "See sections 4.1 and 4.2 of Rosenberg et al. (2012). for details." ;
  		dia_width_err:units = "um" ;
  		dia_width_err:_FillValue = -9999.f ;

  // group attributes:
  		:title = "Size bin calibration of PCASP" ;
  		:comment = "Group containing calibration of size bins of the PCASP. Photodetector voltage pulse-heights are calibrated to the calculated scattering cross-section of known PSL and DEHS monodisperse distributions. Data contained in this group is copied straight from the existing csv calibration files." ;
  		:references = "P.D. Rosenberg, A.R. Dean, P.I. Williams, J.R. Dorsey, A. Minikin, M.A. Pickering and A. Petzold, Particle sizing calibration with refractive index correction for light scattering optical particle counters and impacts upon PCASP and CDP data collected during the Fennec campaign, Atmos. Meas. Tech., 5, 1147-1163, doi:10.5194/amt-5-1147-2012, 2012." ;
  data:

   time = 19082, 19208 ;

   bin = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
      20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30 ;

   applies_to = "C178-C212", "C178-C212" ;

   descr = "ACRUISE-1. MOYA Arctic wetlands. ACSIS-5. ARNA-1", 
      "ACRUISE-1. MOYA Arctic wetlands. ACSIS-5. ARNA-1" ;

   traceability = 
      "269nm (#166237). 303nm (#196947). 345nm (#199283). 400nm (#164245). 453nm (#166631). 508nm (#44115). 600nm (#166837). 707nm (#44582). 799nm (#164766). 903nm (#44869). 0.994um (#200992). 1.101um (#43973). 1.361um (#199629). 1.592um (#204268). 1.745um (#205235). 2.020um (#181058). 2.504um (#190272). 3.007um (#185943).", 
      "269nm (#166237). 303nm (#196947). 345nm (#199283). 400nm (#164245). 453nm (#166631). 508nm (#44115). 600nm (#166837). 707nm (#44582). 799nm (#164766). 903nm (#44869). 0.994um (#200992). 1.101um (#43973). 1.361um (#199629). 1.592um (#204268). 1.745um (#205235). 2.020um (#181058). 2.504um (#190272). 3.007um (#185943)." ;

   cal_flag = 1, 1 ;

   ADC_thres =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

   x-section =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0.450929,
  0.450929, 0.726398,
  0.726398, 0.960547,
  0.960547, 1.64096,
  1.64096, 2.23046,
  2.23046, 2.81721,
  2.81721, 3.41773,
  3.41773, 3.85848,
  3.85848, 4.55542,
  4.55542, 5.25787,
  5.25787, 6.30465,
  6.30465, 7.43958,
  7.43958, 8.6792,
  8.6792, 9.883,
  9.883, 11.3402,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0.0029679,
  0.0029679, 0.00385074,
  0.00385074, 0.00500521,
  0.00500521, 0.00649923,
  0.00649923, 0.0107776,
  0.0107776, 0.017297,
  0.017297, 0.0269402,
  0.0269402, 0.0407034,
  0.0407034, 0.0598088,
  0.0598088, 0.0935149,
  0.0935149, 0.360251,
  0.360251, 0.545627,
  0.545627, 0.703197,
  0.703197, 1.16108,
  1.16108, 1.55778,
  1.55778, 1.95263,
  1.95263, 2.35675,
  2.35675, 2.65336,
  2.65336, 3.12236,
  3.12236, 3.59507,
  3.59507, 4.2995,
  4.2995, 5.06325,
  5.06325, 5.89744,
  5.89744, 6.70754,
  6.70754, 7.68818 ;

   x-section_err =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0,
  0, 0.00703062,
  0.00703062, 0.0155078,
  0.0155078, 0.0381872,
  0.0381872, 0.0575363,
  0.0575363, 0.0767384,
  0.0767384, 0.0963682,
  0.0963682, 0.110768,
  0.110768, 0.133529,
  0.133529, 0.156465,
  0.156465, 0.190636,
  0.190636, 0.227681,
  0.227681, 0.268139,
  0.268139, 0.307426,
  0.307426, 0.354982,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0.000137067,
  0.000137067, 0.000133914,
  0.000133914, 0.000130805,
  0.000130805, 0.000128608,
  0.000128608, 0.000134149,
  0.000134149, 0.000170348,
  0.000170348, 0.000254588,
  0.000254588, 0.000395214,
  0.000395214, 0.000601313,
  0.000601313, 0.000972904,
  0.000972904, 0.0209624,
  0.0209624, 0.0196167,
  0.0196167, 0.0194257,
  0.0194257, 0.0236399,
  0.0236399, 0.0309919,
  0.0309919, 0.0398196,
  0.0398196, 0.0495798,
  0.0495798, 0.0569947,
  0.0569947, 0.0689699,
  0.0689699, 0.0812289,
  0.0812289, 0.0996988,
  0.0996988, 0.119881,
  0.119881, 0.14203,
  0.14203, 0.163605,
  0.163605, 0.189776 ;

   x-section_width =
  -9999, -9999, -9999, -9999, -9999, -9999, -9999, -9999, -9999, -9999, 
      -9999, -9999, -9999, -9999, -9999, -9999, 0.275469, 0.234149, 0.680409, 
      0.589504, 0.58675, 0.600523, 0.440751, 0.696937, 0.702447, 1.04678, 
      1.13493, 1.23961, 1.2038, 1.45723,
  -9999, -9999, -9999, -9999, -9999, -9999, 0.000882833, 0.00115447, 
      0.00149403, 0.00427835, 0.00651938, 0.00964326, 0.0137631, 0.0191054, 
      0.0337061, 0.266736, 0.185376, 0.15757, 0.457879, 0.396705, 0.394852, 
      0.40412, 0.296602, 0.469002, 0.47271, 0.70443, 0.76375, 0.834193, 
      0.810094, 0.980641 ;

   x-section_width_err =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.00898871, 0.00764041, 
      0.0222021, 0.0192358, 0.019146, 0.0195954, 0.0143819, 0.0227414, 
      0.0229212, 0.0341571, 0.0370335, 0.0404492, 0.0392807, 0.0475503,
  _, _, _, _, _, _, 9.87289e-06, 1.29107e-05, 1.6708e-05, 4.78456e-05, 
      7.29075e-05, 0.000107842, 0.000153916, 0.00021366, 0.000376942, 
      0.0071177, 0.00497741, 0.0042308, 0.0122942, 0.0106517, 0.0106019, 
      0.0108508, 0.00796386, 0.0125929, 0.0126924, 0.0189142, 0.0205069, 
      0.0223984, 0.0217513, 0.0263305 ;

   dia_centre =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.591874, 0.729914, 
      0.938788, 1.34543, 1.73936, 1.95487, 2.02668, 2.23672, 2.42188, 
      2.65251, 2.95691, 3.25946, _, _,
  0, 0, 0, 0, 0, 0, 0.164496, 0.17204, 0.180024, 0.192814, 0.210777, 
      0.230073, 0.25094, 0.273276, 0.299024, 0.394132, 0.520465, 0.611762, 
      0.783025, 0.990889, 1.25383, 1.49448, 1.75573, 1.85423, 2.0145, 
      2.17242, 2.36007, 2.57308, 2.76148, 3.05446 ;

   dia_centre_err =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00161694, 0.00366449, 
      0.00404433, 0.0174142, 0.0286537, 0.0267198, 0.0377582, 0.0297179, 
      0.0379129, 0.0465396, 0.080307, 0.05807, _, _,
  0, 0, 0, 0, 0, 0, 0.000669252, 0.000501786, 0.000374634, 0.000267259, 
      0.000260592, 0.000345078, 0.000452744, 0.000554664, 0.000452017, 
      0.00667331, 0.0039655, 0.00127977, 0.00251333, 0.00446769, 0.0265541, 
      0.0277948, 0.0296127, 0.033018, 0.00832448, 0.0177613, 0.032053, 
      0.027667, 0.0255453, 0.0454228 ;

   dia_width =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.151598, 0.124481, 
      0.293265, 0.478078, 0.307111, 0.216725, 0.0740111, 0.159157, 0.181277, 
      0.288284, 0.297718, 0.370406, 0.281908, 0.206015,
  0, 0, 0, 0, 0, 0, 0.00731525, 0.00777243, 0.0081962, 0.017384, 0.0185429, 
      0.0200482, 0.0216851, 0.0229881, 0.0285085, 0.161707, 0.0882481, 
      0.0943458, 0.248179, 0.16755, 0.26987, 0.302136, 0.136449, 0.188126, 
      0.147882, 0.158893, 0.16331, 0.240932, 0.18003, 0.320907 ;

   dia_width_err =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00344668, 0.000662026, 
      0.000364428, 0.0285365, 0.0135932, 0.0139829, 0.0116778, 0.00853104, 
      0.0221077, 0.00964283, 0.042126, 0.0299399, 0.0135907, 0.0468136,
  0, 0, 0, 0, 0, 0, 0.000198556, 0.000163383, 0.000136567, 0.000207127, 
      0.000155022, 0.000132795, 0.000123279, 9.82858e-05, 0.000904034, 
      0.0133466, 0.00228647, 0.00312676, 0.00446463, 0.000615445, 0.0364292, 
      0.0143763, 0.00698934, 0.00989404, 0.0215446, 0.00544942, 0.0209264, 
      0.0138259, 0.0134272, 0.0478624 ;
  } // group bin_cal

group: flow_cal {
  dimensions:
  	time = UNLIMITED ; // (1 currently)
  	max_flows = 256 ;
  variables:
  	float time(time) ;
  		time:standard_name = "time" ;
  		time:long_name = "time of calibration" ;
  		time:timezone = "UTC" ;
  		time:units = "days since 1970-01-01 00:00:00" ;
  		time:strftime_format = "days since %Y-%m-%d %Z" ;
  	string applies_to(time) ;
  		applies_to:long_name = "Each calibration applies to these measurements" ;
  		applies_to:comments = "String of applicable flight numbers for calibration" ;
  	string descr(time) ;
  		descr:long_name = "Description of calibration" ;
  		descr:comment = "Campaign name/s for which these calibrations apply" ;
  	string traceability(time) ;
  		traceability:long_name = "Traceability trail for each calibration" ;
  		traceability:comment = "Calibration of low flow cell s/n 1702010-L" ;
  	int cal_flag(time) ;
  		cal_flag:long_name = "Flag denoting quality of calibration" ;
  		cal_flag:valid_range = 0, 3 ;
  		cal_flag:flag_values = 0, 1, 2, 3 ;
  		cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
  		cal_flag:_FillValue = 3 ;
  	float flows_reported(time, max_flows) ;
  		flows_reported:long_name = "Array of flow rates reported by PCASP for each value in flows_actual" ;
  		flows_reported:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_reported for each time is the same as flows_actual for that time." ;
  		flows_reported:units = "cc/s" ;
  		flows_reported:_FillValue = NaNf ;
  	float flows_actual(time, max_flows) ;
  		flows_actual:long_name = "Array of actual flow rates for each value in flows_reported" ;
  		flows_actual:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_actual for each time is the same as flows_reported for that time." ;
  		flows_actual:units = "cc/s" ;
  		flows_actual:_FillValue = NaNf ;
  	string flow_fit(time) ;
  		flow_fit:long_name = "Calibration equation of sample flow." ;
  		flow_fit:comment = "String of equation used to convert reported flow to calibrated flow rate. This will involve a fit to the data given for the same time stamp in the flows variable. A string is used for flexibility but may be changed to polynomial values in the future if appropriate." ;
  		string flow_fit:_FillValue = "" ;

  // group attributes:
  		:title = "Flow calibration of PCASP" ;
  		:comment = "Gilibrator 2 small cell (to 250cc/m) connected to outlet of PCASP1. Small CV needle valve used to throttle inlet flow with inline Alicat flowmeter used to measure T & P of inlet air" ;
  		:references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
  data:

   time = 17662 ;

   applies_to = "C175-" ;

   descr = _ ;

   traceability = 
      "Calibrated 20170210. Uncertainty of flow = 0.44% + instrument resolution." ;

   cal_flag = 0 ;

   flows_reported =
  1.046, 0.996, 0.911, 0.789, 0.72, 0.611, 0.522, 0.397, 0.334, 0.235, 
      0.148, 0.115, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _ ;

   flows_actual =
  0.919, 0.879, 0.808, 0.699, 0.64, 0.542, 0.455, 0.344, 0.275, 0.185, 
      0.071, 0.022, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _ ;

   flow_fit = "0.280*x**3 - 0.672*x**2 + 1.397*x - 0.123" ;
  } // group flow_cal
}
