netcdf PCASP1_template_calnc {

// This cdl file contains the attributes, dimensions, and variables that are
// applied to all calibration netCDF files for a particular instrument.
//
// This CDL file contains `template` PCASP-1 calibration. Groups for OPAC mixtures
// modified to ignore nucleation and coarse mode particles. RI based on number
// concentration mixture ratios at 80% RH;
//      ACRT. RI = 1.680-3.496e-01i
//      COCL. RI = 1.397-2.328e-03i
//      COAV. RI = 1.589-2.370e-01i
//      COPO. RI = 1.639-2.991e-01i
//      URBA. RI = 1.687-3.583e-01i
//      DESE. RI = 1.399-2.361e-03i
//      MACL. RI = 1.396-2.297e-03i
//      MAPO. RI = 1.600-2.514e-01i
//
// Instrument: PCASP-1
//
// Structure of the cal-nc file is as follows ;
// Global attributes
//  Group: bin_cal
//      Contains scattering cross-section calibration info for size bins.
//    Group: Secondary material sub-group
//      This sub-group of bin_cal/ contains diameter-related variables for
//      another material. Dimensions are inherited from bin_cal. Material
//      information is included in group and variable attributes.
//    Group: Another material sub-group
//      Any number of material sub-groups can be included for different
//      particle types/materials.
//
// author = G. Nott
// email = graeme.nott@faam.ac.uk
// creation = Apr 2023

// global attributes:

    // Universal global file attributes. Do not modify.
    :Conventions = "CF-1.9 ACDD-1.3" ;
    :title = "FAAM calibration data for the PCASP" ;
    :summary = "Bin size and sample flow calibrations for the PCASP relevant to this project." ;
    :instrument = "PCASP-1" ;
    :instrument_model = "Passive Cavity Spectrometer Probe. SPP200 electronics package" ;
    :instrument_manufacturer = "Droplet Measurement Technologies" ;
    :instrument_serial_number = "17884-0190-04" ;
    :references = "https://old.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
//
    :project = "" ;
//
    :source = "Laboratory-based calibration" ;
    :institution = "FAAM Airborne Laboratory" ;
    :creator_institution = "FAAM Airborne Laboratory" ;
    :creator_address = "Building 146, Cranfield University, College Road, Cranfield, Bedford MK43 0AL, UK" ;
    :creator_type = "person" ;
    :creator_name = "Graeme Nott" ;
    :creator_email = "graeme.nott@faam.ac.uk" ;
//    :date_created = "2022-02-10T14:00:00Z" ;
    :publisher_institution = "CEDA" ;
    :publisher_email = "support@ceda.ac.uk" ;
    :publisher_type = "institution" ;
    :publisher_url = "https://www.ceda.ac.uk" ;

    :naming_authority = "uk.ac.faam" ;
//  :id = ;
//  :uuid = ;

//    :revision_date = "2022-02-10T14:00:00Z" ;
    :revision_number = 1 ;
//    :history = "2022-02-10T14:00:00Z cal_ncgen.py v1.0" ;

// ------------------------------------------------------------------------------------
group: bin_cal {
    // Group containing calibration of size bins of the PCASP

    :title = "Size bin calibration of PCASP" ;
    :comment = "Group containing calibration of size bins of the PCASP. Photodetector voltage pulse-heights are calibrated to the calculated scattering cross-section of known PSL and DEHS monodisperse distributions. If one knows the particle refractive index then use the scattering cross-sections for each bin to calculate the bin diameters. For convenience some pre-calculated diameters may be provided in descendant groups, see the group comments for details, although these are intended for quick-look data analysis only. The inclusion of a diameter group does not signify that it is necessarily applicable to any given dataset." ;
    :references = "P.D. Rosenberg, A.R. Dean, P.I. Williams, J.R. Dorsey, A. Minikin, M.A. Pickering and A. Petzold, Particle sizing calibration with refractive index correction for light scattering optical particle counters and impacts upon PCASP and CDP data collected during the Fennec campaign, Atmos. Meas. Tech., 5, 1147-1163, doi:10.5194/amt-5-1147-2012, 2012." ;
    :instrument_collection_angles = "35-120, 60-145 deg" ;
    :instrument_wavelength = "632.8 nm" ;
    :applied = "False" ;

    // Define dimensions for group.
    dimensions:
        time = UNLIMITED ;
        bin = 30 ;
        bin_bounds = 2 ;
        num_gainstages = 3 ;
        polyfit_order = 2 ;

    // Define group coordinate variable
    variables:
        float time(time) ;
            // The units of time may be one of days ('d'), hours ('hr', 'h'),
            // minutes ('min'), or seconds ('sec', 's'). The most appropriate
            // unit given the frequency of calibration should be used.
            time:standard_name = "time" ;
            time:long_name = "time of calibration" ;
            time:units = "days since 1970-01-01 00:00:00 +0000" ;
            time:coverage_content_type = "coordinate" ;
            time:comment = "Multiple calibrations, usually before and after a campaign, may be carried out. A significant difference between the calibrations indicates an instrument alignment change during the campaign. Flag values may indicate a better or worse calibration to apply or else an average of the calibrations could be used." ;

        short bin(bin) ;
            bin:long_name = "bin number" ;
            bin:comment = "The PCASP has 30 bins however the first has a somewhat undefined lower boundary and should therefore usually be discarded." ;
            bin:coverage_content_type = "coordinate" ;

    // Define group variables
        string applies_to(time) ;
            applies_to:long_name = "Calibration applies to this data" ;
            applies_to:comment = "String of applicable flight numbers, dates, or other unique identifier for data that calibration applies to." ;

        string traceability(time) ;
            traceability:long_name = "Traceability of calibration" ;
            traceability:comment = "Information or link to file/s showing traceability of calibration materials and instruments or unique lot numbers for each calibration PSL." ;

        string calibration_file(time) ;
            calibration_file:long_name = "File from which this calibration data has been read" ;

        string source_file(time) ;
            source_file:long_name = "Source file used in calibration processing" ;

        short calibration_qc(time) ;
            calibration_qc:long_name = "Flag denoting quality of calibration" ;
            calibration_qc:valid_range = 0, 3 ;
            calibration_qc:flag_values = 0, 1, 2, 3 ;
            calibration_qc:flag_meanings = "good questionable poor missing_or_bad" ;
            calibration_qc:coverage_content_type = "qualityInformation" ;

        short ADC_threshold(time,bin,bin_bounds) ;
            ADC_threshold:long_name = "Lower and upper analogue-to-digital converter (ADC) thresholds for each bin" ;
            ADC_threshold:comment = "Coverage of each bin in terms of the digitized peak photovoltage. This variable has been included primarily for error checking as the same values should be in the standard data files." ;
            ADC_threshold:valid_range = 0, 12288 ;
            ADC_threshold:coverage_content_type = "auxillaryInformation" ;

        short ADC_range(time,num_gainstages,bin_bounds) ;
            ADC_range:long_name = "Range of analogue-to-digital converter (ADC) values covered by each gain stage" ;
            ADC_range:comment = "Minimum and maximum of ADC values for each gain stage which can be used with corresponding fitting parameters to calculate the scattering cross-section fits for each gain stage" ;
            ADC_range:valid_range = 0, 12288 ;
            ADC_range:coverage_content_type = "auxillaryInformation" ;
            
        float scattering_cross_section(time,bin,bin_bounds) ;
            scattering_cross_section:long_name = "Lower and upper scattering cross-section boundaries for each bin" ;
            scattering_cross_section:comment = "Lower boundary of first bin is undefined." ;
            scattering_cross_section:units = "um**2" ;
            scattering_cross_section:ancillary_variables = "scattering_cross_section_err" ;
            scattering_cross_section:coverage_content_type = "physicalMeasurement" ;

        float scattering_cross_section_err(time,bin,bin_bounds) ;
            scattering_cross_section_err:long_name = "Uncertainty of scattering cross-section boundaries for each bin" ;
            scattering_cross_section_err:comment = "Uncertainties are derived from the uncertainty in the calculated scattering cross-section and the width of the modal bin for each calibration particle. These are discussed in sections 2.1 and 2.23 in Rosenberg et al. [2012] (full citation given in references attribute of this group)." ;
            scattering_cross_section_err:units = "um**2" ;
            scattering_cross_section_err:ancillary_variables = "dependant_scattering_cross_section_err" ;

        float scattering_cross_section_width(time,bin) ;
            scattering_cross_section_width:long_name = "Width of each bin in terms of scattering cross-section" ;
            scattering_cross_section_width:units = "um**2" ;
            scattering_cross_section_width:ancillary_variables = "scattering_cross_section_width_err" ;
            scattering_cross_section_width:coverage_content_type = "physicalMeasurement" ;

        float scattering_cross_section_width_err(time,bin) ;
            scattering_cross_section_width_err:long_name = "Uncertainty of scattering cross-section width for each bin" ;
            scattering_cross_section_width_err:comment = "Uncertainties are derived from the uncertainty in the calculated scattering cross-section and the width of the modal bin for each calibration particle. These are discussed in sections 2.1 and 2.23 in Rosenberg et al. [2012] (full citation given in references attribute of this group)." ;
            scattering_cross_section_width_err:units = "um**2" ;

        short dependant_scattering_cross_section_err(time,bin) ;
            dependant_boundaries:long_name = "Boolean indicator of lower and upper scattering cross-section bin boundary uncertainties being independant/dependant" ;
            dependant_boundaries:comment = "If True (1) then scattering cross-section bin boundary uncertainties are correlated" ;
            dependant_boundaries:valid_range = 0, 1 ;

        float polynomial_fit_parameters(time, num_gainstages,polyfit_order) ;
            polynomial_fit_parameters:long_name = "Polynomial fit parameters of increasing order (eg linear fit is p[0] + p[1]*x) for fitting scattering cross-section to ADC_threshold" ;
            polynomial_fit_parameters:comment = "The PCASP has three gain stages, there is a fit for each gain stage." ;
            polynomial_fit_parameters:ancillary_variables = "polynomial_fit_variance polynomial_fit_covariance" ;

        float polynomial_fit_variance(time,num_gainstages,polyfit_order) ;
            polynomial_fit_variance:long_name = "Variance of each of the polynomial fit parameters" ;

        float polynomial_fit_covariance(time,num_gainstages) ;
            polynomial_fit_covariance:long_name = "Covariance between the polynomial fit parameters" ;


    data:
        // Data is comma-delineated with no additional deliniation between
        // dimensions. Thus the data is presented flattened with the overall
        // length being d1*d2*..dn. As specified in the variable definition,
        // the dimensions are cycled over in reverse order so for multi-
        // dimensional arrays, the last dimension varies fastest. Thus,
        // row-order rather than column order is used for matrices. If
        // var = np.array([[11,12,13],[21,22,23]]) then var.flatten() or
        // np.ravel(var) will write the array in the correct way.
        // Missing data can be written as '_'

        bin = 1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30 ;

//  --------------------------------------------------
    group: ARCT {
        // Group containing calibration of size bins of the PCASP for ARCT aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Arctic (ARCT) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Arctic (ARCT) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.680-3.496e-01i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - ARCT" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.680-3.496e-01i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - ARCT" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.680-3.496e-01i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/ARCT

//  --------------------------------------------------
    group: COCL {
        // Group containing calibration of size bins of the PCASP for COCL aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Continental Clean (COCL) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Continental Clean (COCL) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.397-2.328e-03i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - COCL" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.397-2.328e-03i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - COCL" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.397-2.328e-03i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/COCL

//  --------------------------------------------------
    group: COAV {
        // Group containing calibration of size bins of the PCASP for COAV aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Continental Average (COAV) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Continental Average (COAV) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.589-2.370e-01i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - COAV" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.589-2.370e-01i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - COAV" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.589-2.370e-01i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/COAV


//  --------------------------------------------------
    group: COPO {
        // Group containing calibration of size bins of the PCASP for COPO aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Continental Polluted (COPO) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Continental Polluted (COPO) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.639-2.991e-01i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - COPO" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.639-2.991e-01i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - COPO" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.639-2.991e-01i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/COPO


//  --------------------------------------------------
    group: DESE {
        // Group containing calibration of size bins of the PCASP for DESE aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Desert (DESE) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Desert (DESE) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.399-2.361e-03i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - DESE" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.399-2.361e-03i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - DESE" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.399-2.361e-03i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/DESE


//  --------------------------------------------------
    group: MACL {
        // Group containing calibration of size bins of the PCASP for MACL aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Maritime Clean (MACL) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Maritime Clean (MACL) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.396-2.297e-03i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - MACL" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.396-2.297e-03i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - MACL" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.396-2.297e-03i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/MACL


//  --------------------------------------------------
    group: MAPO {
        // Group containing calibration of size bins of the PCASP for MAPO aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Maritime Polluted (MAPO) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Maritime Polluted (MAPO) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.600-2.514e-01i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - MAPO" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.600-2.514e-01i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - MAPO" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.600-2.514e-01i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/MAPO


//  --------------------------------------------------
    group: URBA {
        // Group containing calibration of size bins of the PCASP for URBA aerosol mix

        :title = "Size bin diameter calibrations based on OPAC Urban (URBA) aerosol mixture. Relative humidity = 0.8." ;
        :comment = "Refractive index for calculation of diameter from scattering cross-section based on the OPAC Urban (URBA) aerosol mixture. Complex refractive indices of the individual aerosol components for 0.65 um (the wavelength in the OPAC tables closest to the PCASP HeNe laser, 0.633 um) were averaged after weighting by the number concentration mixture ratios. Aerosols crudely outside the size range of the instrument are discarded, eg nucleation and coarse mode aerosols, with mixture ratios recalculated before averaging. Spherical particles have been assumed and Mie theory used for the conversion. A relative humidity of 80% has been assumed for water soluble components.\nThis procedure is up for debate, any suggestions or comments please contact the creator. The diameter size bin boundaries are intended for quick-look data only, it remains up to the user to decide if it is suitable for their particular scenario. Feel free to contact the creator to discuss applicability.\n\nRefractive index = 1.687-3.583e-01i." ;
        :references = "https://geisa.aeris-data.fr/opac/. Hess, M., Koepke, P., & Schult, I. (1998). Optical Properties of Aerosols and Clouds: The Software Package OPAC, Bulletin of the American Meteorological Society, 79(5), 831-844, doi:10.1175/1520-0477(1998)079<0831:OPOAAC>2.0.CO;2." ;

        // Define group variables
        variables:

            string calibration_file(time) ;
                calibration_file:long_name = "File from which this calibration data has been read" ;

            string source_file(time) ;
                source_file:long_name = "Source file used in calibration processing" ;

            float diameter_centre(time,bin) ;
                diameter_centre:long_name = "Centre diameter of each bin for given aerosol mixture - URBA" ;
                diameter_centre:comment = "Weighted average of all diameter region centres covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_centre:refractive_index = "1.687-3.583e-01i" ;
                diameter_centre:shape = "spherical" ;
                diameter_centre:units = "um" ;
                diameter_centre:ancillary_variables = "diameter_centre_err dia_width" ;
                diameter_centre:coverage_content_type = "physicalMeasurement" ;

            float diameter_centre_err(time,bin) ;
                diameter_centre_err:long_name = "Uncertainty of bin centre diameter" ;
                diameter_centre_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_centre_err:units = "um" ;
                diameter_centre_err:coverage_content_type = "physicalMeasurement" ;

            float diameter_width(time,bin) ;
                diameter_width:long_name = "Width in terms of diameter of each bin for given aerosol mixture - URBA" ;
                diameter_width:comment = "Sum of all diameter regions covered by the scattering cross-sections of each bin. This is discussed in sections 4.1 and 4.2 in Rosenberg et al. [2012]" ;
                diameter_width:refractive_index = "1.687-3.583e-01i" ;
                diameter_width:shape = "spherical" ;
                diameter_width:units = "um" ;
                diameter_width:ancillary_variables = "diameter_width_err" ;
                diameter_width:coverage_content_type = "physicalMeasurement" ;

            float diameter_width_err(time,bin) ;
                diameter_width_err:long_name = "Uncertainty of bin diameter width" ;
                diameter_width_err:comment = "Uncertainties are discussed in sections 4.1 and 4.2 in Rosenberg et al." ;
                diameter_width_err:units = "um" ;
                diameter_width_err:coverage_content_type = "physicalMeasurement" ;

        } // End group bin_cal/URBA

    } // End group bin_cal



// ------------------------------------------------------------------------------------
group: flow_cal {
    // Group containing calibration of flow rates of the PCASP
    //
    :title = "Sample flow calibration of PCASP" ;
    :comment = "The PCASP sample flow was choked by an Alicat MC flow controller with a Gilibrator 3 dry cell flow calibrator connected to the outlet of the PCASP sample flow meter. Volumetric flow (accuracy +/-1%%) was averaged over 10-20 samples over a range of flow rates. Standard condition flows were calculated using the Gilibrator temperature (+/-0.3%%) and pressure (+/-4.5 mbar) sensors and compared with standard flow of PCASP sample flow (Honeywell AWM3100V, +/-0.5%%) as reported by PADS." ;
    :references = "http://old.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
    :applied = "True" ;

    // The units of time may be one of days ('d'), hours ('hr', 'h'),
    // minutes ('min'), or seconds ('sec', 's') and the most appropriate unit
    // for the frequency of calibration should be used.
    dimensions:
        time = UNLIMITED ;
        max_flows = 32 ;    // Maximum number of different flows in a calibration

    // Define group coordinate variable
    variables:
        float time(time) ;
            // The units of time may be one of days ('d'), hours ('hr', 'h'),
            // minutes ('min'), or seconds ('sec', 's') and the most appropriate
            // unit for the frequency of calibration should be used.
            time:standard_name = "time" ;
            time:long_name = "time of calibration" ;
            time:timezone = "UTC" ;
            time:units = "days since 1970-01-01 00:00:00" ;
            time:strftime_format = "days since %Y-%m-%d %H:%M:%S%Z" ;

    // Define group variables
        string applies_to(time) ;
            applies_to:long_name = "Calibration applies to this data" ;
            applies_to:comments = "String of applicable flight numbers, dates, or other unique identifier for data that calibration applies to." ;

        string traceability(time) ;
            traceability:long_name = "Traceability of calibration" ;
            traceability:comment = "Links to calibration certificates or other identifiers showing traceability of calibration instruments." ;

        short calibration_qc(time) ;
            calibration_qc:long_name = "Flag denoting quality of calibration" ;
            calibration_qc:valid_range = 0, 3 ;
            calibration_qc:flag_values = 0, 1, 2, 3 ;
            calibration_qc:flag_meanings = "good questionable poor missing_or_bad" ;
            calibration_qc:_FillValue = 3 ;
            calibration_qc:coverage_content_type = "qualityInformation" ;

        float flows_reported(time,max_flows) ;
            flows_reported:long_name = "Sample flow rate reported by PCASP for each value in flows_actual" ;
            flows_reported:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the length of flows_reported for each time is the same as flows_actual for that time." ;
            flows_reported:units = "scc/s" ;
//            flows_reported:valid_min = -0.01 ;
            flows_reported:_FillValue = -999.9f ;
            flows_reported:coverage_content_type = "physicalMeasurement" ;

        float flows_actual(time,max_flows) ;
            flows_actual:long_name = "Verified sample flow rate for each value in flows_reported" ;
            flows_actual:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_actual for each time is the same as flows_reported for that time." ;
            flows_actual:units = "scc/s" ;
//            flows_actual:valid_min = -0.01 ;
            flows_actual:_FillValue = -999.9f ;
            flows_actual:coverage_content_type = "physicalMeasurement" ;

        string flow_fit(time) ;
            flow_fit:long_name = "Calibration equation of sample flow" ;
            flow_fit:comment = "String of equation used to convert reported sample flow to calibrated sample flow rate. It is assumed that the same conversion can be used for standard conditions and volumetric flows." ;
            flow_fit:_FillValue = "" ;


    data:
        // Data is comma-delineated with no additional deliniation between
        // dimensions. Thus the data is presented flattened with the overall
        // length being d1*d2*..dn. As specified in the variable definition,
        // the dimensions are cycled over in reverse order so for multi-
        // dimensional arrays, the last dimension varies fastest. Thus,
        // row-order rather than column order is used for matrices.. If
        // var = np.array([[11,12,13],[21,22,23]]) then var.flatten() or
        // np.ravel(var) will write the array in the correct way.

    } // End group flow_cal

} // EOF
