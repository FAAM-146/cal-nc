netcdf PCASP_faam_20191107_v001_r000_cal {

// global attributes:
		:Conventions = "CF-1.6" ;
		:institution = "FAAM. Facility for Airborne Atmospheric Measurements" ;
		:address = "Building 146, Cranfield University, Cranfield MK43 0AL UK" ;
		:title = "FAAM calibration data for the PCASP-2" ;
		:source = "Laboratory-based calibration" ;
		:instr = "PCASP-2" ;
		:instr_long_name = "Passive Cavity Spectrometer Probe. SPP200 electronics package" ;
		:instr_serialnumber = "PMI-1022-1202-31" ;
		:references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
		:username = "Graeme Nott <graeme.nott@faam.ac.uk>" ;
		:history = "20191202T1747 Initial creation" ;
		:software_version = "0.3" ;

group: bin_cal {
  dimensions:
  	time = UNLIMITED ; // (2 currently)
  	bin = 30 ;
  	bin_bounds = 2 ;
  variables:
  	float time(time) ;
  		time:standard_name = "time" ;
  		time:long_name = "time of calibration" ;
  		time:timezone = "UTC" ;
  		time:units = "days since 1970-01-01 00:00:00" ;
  		time:strftime_format = "days since %Y-%m-%d %Z" ;
  	int bin(bin) ;
  		bin:long_name = "bin number" ;
  		bin:comment = "The PCASP has 30 bins however the first has a somewhat undefined lower boundary and should therefore be discarded." ;
  	string applies_to(time) ;
  		applies_to:long_name = "Each calibration applies to these measurements" ;
  		applies_to:comment = "String of applicable flight numbers for calibration" ;
  	string descr(time) ;
  		descr:long_name = "Description of calibration" ;
  		descr:comment = "Campaign name/s for which these calibrations apply" ;
  	string traceability(time) ;
  		traceability:long_name = "Traceability trail for each calibration" ;
  		traceability:comment = "Unique lot numbers for each calibration PSL. These can be traced to the original NIST-traceable certificates." ;
  	int cal_flag(time) ;
  		cal_flag:long_name = "Flag denoting quality of calibration" ;
  		cal_flag:valid_range = 0, 3 ;
  		cal_flag:flag_values = 0, 1, 2, 3 ;
  		cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
  		cal_flag:_FillValue = 3 ;
  	int ADC_thres(time, bin, bin_bounds) ;
  		ADC_thres:long_name = "Lower and upper ADC thresholds for each bin" ;
  		ADC_thres:comment = "Coverage of each bin in terms of the digitized peak photovoltage. This variable has been included primarily for error checking as the same values should be in the standard data files." ;
  		ADC_thres:valid_range = 0, 1288 ;
  		ADC_thres:_FillValue = -2147483648 ;
  	float x-section(time, bin, bin_bounds) ;
  		x-section:long_name = "Scattering cross-section boundaries for each bin" ;
  		x-section:comment = "Lower boundary of first bin is undefined." ;
  		x-section:units = "m**2" ;
  		x-section:ancillary_variables = "x-section_width_err" ;
  		x-section:_FillValue = -9999.f ;
  	float x-section_err(time, bin, bin_bounds) ;
  		x-section_err:long_name = "Uncertainty of scattering cross section boundaries for each bin" ;
  		x-section_err:comment = "Straight-line fits for scattering cross-section versus ADC voltage are calculated along with sensitivities to the uncertainty in these data. See section 2.2.3 of Rosenberg et al. (2012) for details." ;
  		x-section_err:_FillValue = -9999.f ;
  	float x-section_width(time, bin) ;
  		x-section_width:long_name = "Width of each bin in terms of scattering cross section" ;
  	float x-section_width_err(time, bin) ;
  		x-section_width_err:long_name = "Uncertainty of scattering cross section boundaries for each bin" ;
  		x-section_width_err:comment = "" ;
  		x-section_width_err:flag_values = 0, 1 ;
  		x-section_width_err:flag_meanings = "Independent_uncertainties \n                                             Dependent_uncertainties" ;
  		x-section_width_err:_FillValue = -9999.f ;
  	float dia_centre(time, bin) ;
  		dia_centre:long_name = "Centre diameter associated with each bin number for given particle material properties" ;
  		dia_centre:comment = "This is the weighted average of each of the regions of the scattering curve which include the range of scattering cross-sections in each bin with the uncertainty of these boundaries included. This is discussed in sections 4.1 and 4.2 of Rosenberg et al. (2012)." ;
  		dia_centre:refractive_index = "1.59+0i" ;
  		dia_centre:shape = "spherical" ;
  		dia_centre:units = "um" ;
  		dia_centre:ancillary_variables = "dia_centre_err dia_width" ;
  		dia_centre:_FillValue = -9999.f ;
  	float dia_centre_err(time, bin) ;
  		dia_centre_err:long_name = "Uncertainty of bin centre diameter" ;
  		dia_centre_err:comment = "See sections 4.1 and 4.2 of Rosenberg et al. (2012). for details." ;
  		dia_centre_err:units = "um" ;
  		dia_centre_err:_FillValue = -9999.f ;
  	float dia_width(time, bin) ;
  		dia_width:long_name = "Diameter width associated with each bin number for given particle material properties" ;
  		dia_width:comment = "This is the sum of all regions of the scattering curve which include the range of scattering cross-sections in each bin with the uncertainty of these boundaries included. This is discussed in sections 4.1 and 4.2 of Rosenberg et al. (2012)." ;
  		dia_width:refractive_index = "1.59+0i" ;
  		dia_width:shape = "spherical" ;
  		dia_width:units = "um" ;
  		dia_width:ancillary_variables = "dia_width_err" ;
  		dia_width:_FillValue = -9999.f ;
  	float dia_width_err(time, bin) ;
  		dia_width_err:long_name = "Uncertainty of bin width" ;
  		dia_width_err:comment = "See sections 4.1 and 4.2 of Rosenberg et al. (2012). for details." ;
  		dia_width_err:units = "um" ;
  		dia_width_err:_FillValue = -9999.f ;

  // group attributes:
  		:title = "Size bin calibration of PCASP" ;
  		:comment = "Group containing calibration of size bins of the PCASP. Photodetector voltage pulse-heights are calibrated to the calculated scattering cross-section of known PSL and DEHS monodisperse distributions. Data contained in this group is copied straight from the existing csv calibration files." ;
  		:references = "P.D. Rosenberg, A.R. Dean, P.I. Williams, J.R. Dorsey, A. Minikin, M.A. Pickering and A. Petzold, Particle sizing calibration with refractive index correction for light scattering optical particle counters and impacts upon PCASP and CDP data collected during the Fennec campaign, Atmos. Meas. Tech., 5, 1147-1163, doi:10.5194/amt-5-1147-2012, 2012." ;
  data:

   time = 18082, 18208 ;

   bin = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
      20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30 ;

   applies_to = "C178-C212", "C178-C212" ;

   descr = 
      "ACRUISE-1. MOYA Arctic wetlands. ACSIS-5. ARNA-1. DMA u/s. PSLs for mid-gain stage.", 
      "ACRUISE-1. MOYA Arctic wetlands. ACSIS-5. ARNA-1. High-gain stage card u/s. Fine in flight-blew in lab?" ;

   traceability = 
      "125nm (#44245). 150nm (#202026). 203nm (#44793). 216nm (#16779). 240nm (#45059). 269nm (#166237). 303nm (#196947). 345nm (#199283). 400nm (#164245). 453nm (#166631). 508nm (#44115). 600nm (#166837). 707nm (#44582). 799nm (#164766). 903nm (#44869). 0.994um (#200992). 1.101um (#43973). 1.361um (#199629). 1.592um (#204268). 1.745um (#205235). 2.020um (#181058). 2.504um (#190272). 3.007um (#185943).", 
      "269nm (#166237). 303nm (#196947). 345nm (#199283). 400nm (#164245). 453nm (#166631). 508nm (#44115). 600nm (#166837). 707nm (#44582). 799nm (#164766). 903nm (#44869). 0.994um (#200992). 1.101um (#43973). 1.361um (#199629). 1.592um (#204268). 1.745um (#205235). 2.020um (#181058). 2.504um (#190272). 3.007um (#185943)." ;

   cal_flag = 1, 1 ;

   ADC_thres =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

   x-section =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0.00254097,
  0.00254097, 0.00373883,
  0.00373883, 0.00530527,
  0.00530527, 0.00733242,
  0.00733242, 0.0131375,
  0.0131375, 0.0219832,
  0.0219832, 0.0350676,
  0.0350676, 0.053742,
  0.053742, 0.079665,
  0.079665, 0.125399,
  0.125399, 0.485015,
  0.485015, 0.741009,
  0.741009, 0.958605,
  0.958605, 1.59091,
  1.59091, 2.13874,
  2.13874, 2.68401,
  2.68401, 3.24208,
  3.24208, 3.65167,
  3.65167, 4.29933,
  4.29933, 4.95212,
  4.95212, 5.9249,
  5.9249, 6.9796,
  6.9796, 8.13157,
  8.13157, 9.25027,
  9.25027, 10.6045,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0.0029679,
  0.0029679, 0.00385074,
  0.00385074, 0.00500521,
  0.00500521, 0.00649923,
  0.00649923, 0.0107776,
  0.0107776, 0.017297,
  0.017297, 0.0269402,
  0.0269402, 0.0407034,
  0.0407034, 0.0598088,
  0.0598088, 0.0935149,
  0.0935149, 0.360251,
  0.360251, 0.545627,
  0.545627, 0.703197,
  0.703197, 1.16108,
  1.16108, 1.55778,
  1.55778, 1.95263,
  1.95263, 2.35675,
  2.35675, 2.65336,
  2.65336, 3.12236,
  3.12236, 3.59507,
  3.59507, 4.2995,
  4.2995, 5.06325,
  5.06325, 5.89744,
  5.89744, 6.70754,
  6.70754, 7.68818 ;

   x-section_err =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0.000842166,
  0.000842166, 0.000787564,
  0.000787564, 0.000722996,
  0.000722996, 0.00065436,
  0.00065436, 0.000595998,
  0.000595998, 0.000898705,
  0.000898705, 0.00165073,
  0.00165073, 0.00283561,
  0.00283561, 0.00452195,
  0.00452195, 0.00752266,
  0.00752266, 0.012612,
  0.012612, 0.0136605,
  0.0136605, 0.0189594,
  0.0189594, 0.0405093,
  0.0405093, 0.0607357,
  0.0607357, 0.0811873,
  0.0811873, 0.102249,
  0.102249, 0.117751,
  0.117751, 0.142306,
  0.142306, 0.167087,
  0.167087, 0.20405,
  0.20405, 0.244153,
  0.244153, 0.287975,
  0.287975, 0.330541,
  0.330541, 0.38208,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, 0.000137067,
  0.000137067, 0.000133914,
  0.000133914, 0.000130805,
  0.000130805, 0.000128608,
  0.000128608, 0.000134149,
  0.000134149, 0.000170348,
  0.000170348, 0.000254588,
  0.000254588, 0.000395214,
  0.000395214, 0.000601313,
  0.000601313, 0.000972904,
  0.000972904, 0.0209624,
  0.0209624, 0.0196167,
  0.0196167, 0.0194257,
  0.0194257, 0.0236399,
  0.0236399, 0.0309919,
  0.0309919, 0.0398196,
  0.0398196, 0.0495798,
  0.0495798, 0.0569947,
  0.0569947, 0.0689699,
  0.0689699, 0.0812289,
  0.0812289, 0.0996988,
  0.0996988, 0.119881,
  0.119881, 0.14203,
  0.14203, 0.163605,
  0.163605, 0.189776 ;

   x-section_width =
  -9999, -9999, -9999, -9999, -9999, -9999, 0.00119786, 0.00156644, 
      0.00202715, 0.00580503, 0.00884576, 0.0130844, 0.0186744, 0.025923, 
      0.0457338, 0.359616, 0.255995, 0.217595, 0.632307, 0.547828, 0.545268, 
      0.558068, 0.409591, 0.647666, 0.652786, 0.972779, 1.0547, 1.15198, 
      1.1187, 1.35421,
  -9999, -9999, -9999, -9999, -9999, -9999, 0.000882833, 0.00115447, 
      0.00149403, 0.00427835, 0.00651938, 0.00964326, 0.0137631, 0.0191054, 
      0.0337061, 0.266736, 0.185376, 0.15757, 0.457879, 0.396705, 0.394852, 
      0.40412, 0.296602, 0.469002, 0.47271, 0.70443, 0.76375, 0.834193, 
      0.810094, 0.980641 ;

   x-section_width_err =
  _, _, _, _, _, _, 7.89979e-05, 0.000103305, 0.000133689, 0.000382836, 
      0.000583369, 0.0008629, 0.00123156, 0.0017096, 0.0030161, 0.01394, 
      0.00974825, 0.00828601, 0.0240782, 0.0208613, 0.0207638, 0.0212512, 
      0.0155972, 0.0246631, 0.024858, 0.0370434, 0.0401628, 0.0438671, 
      0.0425999, 0.0515682,
  _, _, _, _, _, _, 9.87289e-06, 1.29107e-05, 1.6708e-05, 4.78456e-05, 
      7.29075e-05, 0.000107842, 0.000153916, 0.00021366, 0.000376942, 
      0.0071177, 0.00497741, 0.0042308, 0.0122942, 0.0106517, 0.0106019, 
      0.0108508, 0.00796386, 0.0125929, 0.0126924, 0.0189142, 0.0205069, 
      0.0223984, 0.0217513, 0.0263305 ;

   dia_centre =
  0, 0, 0, 0, 0, 0, 0.161532, 0.172353, 0.182843, 0.198507, 0.219736, 
      0.242032, 0.265824, 0.290497, 0.3175, 0.430883, 0.601522, 0.732623, 
      0.935458, 1.31996, 1.68059, 1.89863, 2.0102, 2.17978, 2.34456, 2.56224, 
      2.80224, 3.14323, _, _,
  0, 0, 0, 0, 0, 0, 0.164496, 0.17204, 0.180024, 0.192814, 0.210777, 
      0.230073, 0.25094, 0.273276, 0.299024, 0.394132, 0.520465, 0.611762, 
      0.783025, 0.990889, 1.25383, 1.49448, 1.75573, 1.85423, 2.0145, 
      2.17242, 2.36007, 2.57308, 2.76148, 3.05446 ;

   dia_centre_err =
  0, 0, 0, 0, 0, 0, 0.00545099, 0.00334094, 0.0019438, 0.00057022, 
      0.000782926, 0.00181591, 0.00268728, 0.0033132, 0.00264808, 0.00329778, 
      0.00056109, 0.00306263, 0.00460748, 0.0181687, 0.0453911, 0.0394052, 
      0.00746736, 0.0348722, 0.0412279, 0.0449035, 0.0693954, 0.0622692, _, _,
  0, 0, 0, 0, 0, 0, 0.000669252, 0.000501786, 0.000374634, 0.000267259, 
      0.000260592, 0.000345078, 0.000452744, 0.000554664, 0.000452017, 
      0.00667331, 0.0039655, 0.00127977, 0.00251333, 0.00446769, 0.0265541, 
      0.0277948, 0.0296127, 0.033018, 0.00832448, 0.0177613, 0.032053, 
      0.027667, 0.0255453, 0.0454228 ;

   dia_width =
  0, 0, 0, 0, 0, 0, 0.0110807, 0.0105606, 0.0104203, 0.0209073, 0.021551, 
      0.0230407, 0.024543, 0.0248039, 0.0292088, 0.197556, 0.144091, 
      0.118111, 0.287558, 0.432708, 0.288753, 0.228328, 0.09849, 0.147777, 
      0.139107, 0.274045, 0.238714, 0.393081, 0.266215, 0.282616,
  0, 0, 0, 0, 0, 0, 0.00731525, 0.00777243, 0.0081962, 0.017384, 0.0185429, 
      0.0200482, 0.0216851, 0.0229881, 0.0285085, 0.161707, 0.0882481, 
      0.0943458, 0.248179, 0.16755, 0.26987, 0.302136, 0.136449, 0.188126, 
      0.147882, 0.158893, 0.16331, 0.240932, 0.18003, 0.320907 ;

   dia_width_err =
  0, 0, 0, 0, 0, 0, 0.00261851, 0.00163823, 0.00116194, 0.00158655, 
      0.00111861, 0.000947636, 0.00079547, 0.00045792, 0.00529615, 
      0.00659557, 0.00406565, 0.000949336, 0.00267623, 0.0324692, 0.0111308, 
      0.00933062, 0.0273542, 0.0117725, 0.019486, 0.0114616, 0.031484, 
      0.0313069, 0.0150962, 0.0280426,
  0, 0, 0, 0, 0, 0, 0.000198556, 0.000163383, 0.000136567, 0.000207127, 
      0.000155022, 0.000132795, 0.000123279, 9.82858e-05, 0.000904034, 
      0.0133466, 0.00228647, 0.00312676, 0.00446463, 0.000615445, 0.0364292, 
      0.0143763, 0.00698934, 0.00989404, 0.0215446, 0.00544942, 0.0209264, 
      0.0138259, 0.0134272, 0.0478624 ;
  } // group bin_cal

group: flow_cal {
  dimensions:
  	time = UNLIMITED ; // (1 currently)
  	max_flows = 64 ;
  variables:
  	float time(time) ;
  		time:standard_name = "time" ;
  		time:long_name = "time of calibration" ;
  		time:timezone = "UTC" ;
  		time:units = "days since 1970-01-01 00:00:00" ;
  		time:strftime_format = "days since %Y-%m-%d %Z" ;
  	string applies_to(time) ;
  		applies_to:long_name = "Each calibration applies to these measurements" ;
  		applies_to:comments = "String of applicable flight numbers for calibration" ;
  	string descr(time) ;
  		descr:long_name = "Description of calibration" ;
  		descr:comment = "Campaign name/s for which these calibrations apply" ;
  	string traceability(time) ;
  		traceability:long_name = "Traceability trail for each calibration" ;
  		traceability:comment = "Calibration of low flow cell s/n 1702010-L" ;
  	int cal_flag(time) ;
  		cal_flag:long_name = "Flag denoting quality of calibration" ;
  		cal_flag:valid_range = 0, 3 ;
  		cal_flag:flag_values = 0, 1, 2, 3 ;
  		cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
  		cal_flag:_FillValue = 3 ;
  	float flows_reported(time, max_flows) ;
  		flows_reported:long_name = "Array of flow rates reported by PCASP for each value in flows_actual" ;
  		flows_reported:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_reported for each time is the same as flows_actual for that time." ;
  		flows_reported:units = "cc/s" ;
  		flows_reported:_FillValue = NaNf ;
  	float flows_actual(time, max_flows) ;
  		flows_actual:long_name = "Array of actual flow rates for each value in flows_reported" ;
  		flows_actual:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_actual for each time is the same as flows_reported for that time." ;
  		flows_actual:units = "cc/s" ;
  		flows_actual:_FillValue = NaNf ;
  	string flow_fit(time) ;
  		flow_fit:long_name = "Calibration equation of sample flow." ;
  		flow_fit:comment = "String of equation used to convert reported flow to calibrated flow rate. This will involve a fit to the data given for the same time stamp in the flows variable. A string is used for flexibility but may be changed to polynomial values in the future if appropriate." ;
  		string flow_fit:_FillValue = "" ;

  // group attributes:
  		:title = "Flow calibration of PCASP" ;
  		:comment = "Gilibrator 2 small cell (to 250cc/m) connected to outlet of PCASP1. Small CV needle valve used to throttle inlet flow with inline Alicat flowmeter used to measure T & P of inlet air" ;
  		:references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
  data:

   time = 17660 ;

   applies_to = "C173-" ;

   descr = _ ;

   traceability = 
      "Calibrated 20170210. Uncertainty of flow = 0.44% + instrument resolution." ;

   cal_flag = 0 ;

   flows_reported =
  1.046, 0.996, 0.911, 0.789, 0.72, 0.611, 0.522, 0.397, 0.334, 0.235, 
      0.148, 0.115, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _ ;

   flows_actual =
  0.919, 0.879, 0.808, 0.699, 0.64, 0.542, 0.455, 0.344, 0.275, 0.185, 
      0.071, 0.022, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _ ;

   flow_fit = "0.280*x**3 - 0.672*x**2 + 1.397*x - 0.123" ;
  } // group flow_cal
}
