netcdf PCASP1_cal_20180117 {

// This cdl file contains the attributes, dimensions, and variables that are
// applied to all calibration netCDF files for a particular instrument. This
// file combined with FAAMheader.cdl provides the source data for PCASP1 
// calibration netCDF files. Some of these fields shall be modified/
// overwritten by cal_ncgen.py if it is used.
//
// author = G. Nott
// email = graeme.nott@faam.ac.uk
// creation = Jan 2018

// global attributes:
    
    // Universal global file attributes. Do not modify.
    :Conventions = "CF-1.6";
    :NCO = "4.1.3";
    :_Format = "netCDF-4";
    :institution = "FAAM. Facility for Airborne Atmospheric Measurements";
    :address = "Building 146, Cranfield University, Cranfield MK43 0AL UK";

    // Instrument global file attributes. 
    :title = "FAAM calibration data for the PCASP-1";
    :source = "Laboratory-based calibration";
    :instr = "PCASP-1";
    :instr_long_name = "Passive Cavity Spectrometer Probe. SPP200 electronics package";
    :instr_serialnumber = "17884-0190-04";
    :references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp";

// The following global attributes shall be modified by cal_ncgen.py if used
    :username = "graeme.nott@faam.ac.uk, Graeme Nott";
    :history = "20180111";

// Define global dimensions for generated file.
// calnc files have a root unlimited dimension of time. The units of time may
// be one of days ('d'), hours ('hr', 'h'), minutes ('min'), or seconds ('sec',
// 's') and the most appropriate unit for the frequency of calibration should
// be used.
dimensions:
    time = UNLIMITED ; // (2 currently)

// Define global coordinate variable
variables:
    float time(time);
    time:standard_name = "time";
    time:long_name = "time of calibration";
    time:timezone = "UTC";
    time:units = "days since 2010-01-01 00:00:00";
    time:strftime_format = "days since %Y-%m-%d %H:%M:%S%Z";

data:
    time = 2818.5, 2864.5;

group: bin_cal {
    // Group containing calibration of size bins of the PCASP
    //
    :title = "Size bin calibration of PCASP";
    :comment = "Group containing calibration of size bins of the PCASP. Photodetector voltage pulse-heights are calibrated to the calculated scattering cross-section of known PSL and DEHS monodisperse distributions.";
    :references = "P.D. Rosenberg, A.R. Dean, P.I. Williams, J.R. Dorsey, A. Minikin, M.A. Pickering and A. Petzold, Particle sizing calibration with refractive index correction for light scattering optical particle counters and impacts upon PCASP and CDP data collected during the Fennec campaign, Atmos. Meas. Tech., 5, 1147-1163, doi:10.5194/amt-5-1147-2012, 2012.";

    // Define any group dimensions in addition to the global dimension, time
    dimensions:
        bin = 30;
        bin_bounds = 2;

    // Define group coordinate variable
    variables:
        int bin(bin);
            bin:long_name = "bin number";

    // Define group variables
        string applies_to(time);
            applies_to:long_name = "Each calibration applies to these measurements";
            applies_to:comments = "String of applicable flight numbers for each calibration date";

        string traceability(time);
            traceability:long_name = "Traceability trail for each calibration";
            traceability:comment = "Link to file/s showing traceability of calibration materials and instruments";

        int cal_flag(time);
            cal_flag:long_name = "Flag denoting quality of calibration";
            cal_flag:valid_range = 0, 3;
            cal_flag:flag_values = 0, 1, 2, 3;
            cal_flag:flag_meanings = "good questionable poor missing_or_bad";
            cal_flag:_FillValue = 3;

        int ADC_thres(time,bin,bin_bounds);
            ADC_thres:long_name = "Lower and upper ADC thresholds for each bin";
            ADC_thres:comment = "Coverage of each bin in terms of the digitized peak photovoltage. This variable has been included primarily for error checking as the same vaules should be in the standard data files.";
            ADC_thres:valid_range = 0, 1288;
            ADC_thres:_FillValue = NaN;

        float x-section(time,bin,bin_bounds);
            x-section:long_name = "Scattering cross-section boundaries for each bin";
            x-section:comment = "Lower boundary of first bin is undefined.";
            x-section:units = "m**2";
            x-section:ancillary_variables = "x-section_err";
            x-section:_FillValue = NaN;

        float x-section_err(time,bin,bin_bounds);
            x-section_err:long_name = "Uncertainty of scattering cross section boundaries for each bin";
            x-section_err:comment = "Comment here about calculation of uncertainties";
            x-section_err:_FillValue = "NaN";

        float x-section_width(time,bin);
            x-section_width:long_name = "Width of each bin in terms of scattering cross section";
            x-section:units = "m**2";
            x-section:ancillary_variables = "x-section_width_err";
            x-section:_FillValue = "NaN";

        float x-section_width_err(time,bin);
            x-section_width_err:long_name = "Uncertainty of scattering cross section boundaries for each bin";
            x-section_width_err:comment = "Comment here about calculation of uncertainties";
            x-section_width_err:flag_values = 0, 1;
            x-section_width_err:flag_meanings = "Independent_uncertainties 
                                                 Dependent_uncertainties";
            x-section_width_err:_FillValue = "NaN";

        float dia_centre(time,bin);
            dia_centre:long_name = "Centre diameter associated with each bin number for given particle material properties";
            dia_centre:comment = "Comments here about the derivation of diameter";
            dia_centre:refractive_index = "1.59+0i";
            dia_centre:shape = "spherical";
            dia_centre:units = "um";
            dia_centre:ancillary_variables = "dia_centre_err dia_width";
            dia_centre:_FillValue = "NaN";

        float dia_centre_err(time,bin);
            dia_centre_err:long_name = "Uncertainty of bin centre diameter";
            dia_centre_err:comment = "Comment here about calculation of uncertainties";
            dia_centre_err:units = "um";
            dia_centre_err:_FillValue = "NaN";

        float dia_width(time,bin);
            dia_width:long_name = "Diameter width associated with each bin number for given particle material properties";
            dia_width:comment = "Comments here about the derivation of diameter";
            dia_width:refractive_index = "1.59+0i";
            dia_width:shape = "spherical";
            dia_width:units = "um";
            dia_width:ancillary_variables = "dia_width_err";
            dia_width:_FillValue = "NaN";

        float dia_width_err(time,bin);
            dia_width_err:long_name = "Uncertainty of bin width";
            dia_width_err:comment = "Comment here about calculation of uncertainties";
            dia_width_err:units = "um";
            dia_width_err:_FillValue = "NaN";


    data:
        // Data is comma-delineated with no additional deliniation between 
        // dimensions. Thus the data is presented flattened with the overall 
        // length being d1*d2*..dn. As specified in the variable definition,
        // the dimensions are cycled over in reverse order so for multi-
        // dimensional arrays, the last dimension varies fastest. Thus, 
        // row-order rather than column order is used for matrices.. If 
        // var = np.array([[11,12,13],[21,22,23]]) then var.flatten() or 
        // np.ravel(var) will write the array in the correct way.
        // Missing data can be written as '_'

        applies_to = "C027-C055", "C057-C071";
        traceability = "","";
        cal_flag = 0, 0;

        ADC_thres = _, 692,692, 1146,1146, 1814,1814, 2769,2769, 4096,4096, 4192,4192, 4231,4231, 4282,4282, 4348,4348, 4537,4537, 4825,4825, 5251,5251, 5859,5859, 6703,6703, 8192,8192, 8335,8335, 8435,8435, 8520,8520, 8767,8767, 8981,8981, 9194,9194, 9412,9412, 9572,9572, 9825,9825, 10080,10080, 10460,10460, 10872,10872, 11322,11322, 11759,11759, 12288,
                            _, 692,692, 1146,1146, 1814,1814, 2769,2769, 4096,4096, 4192,4192, 4231,4231, 4282,4282, 4348,4348, 4537,4537, 4825,4825, 5251,5251, 5859,5859, 6703,6703, 8192,8192, 8335,8335, 8435,8435, 8520,8520, 8767,8767, 8981,8981, 9194,9194, 9412,9412, 9572,9572, 9825,9825, 10080,10080, 10460,10460, 10872,10872, 11322,11322, 11759,11759, 12288 ;

        x-section = _, 0.000484975,
                    0.000484975,0.000582489,
                    0.000582489, 0.000725968,
                    0.000725968, 0.00093101,
                    0.0009311, 0.00121611,
                    0.00121611, 0.00156032,
                    0.00156032, 0.0021721,
                    0.0021721, 0.00297209,
                    0.00297209, 0.00400738,
                    0.00400738, 0.00697209,
                    0.00697209, 0.0114897,
                    0.0114897, 0.0181721,
                    0.0181721, 0.0277093,
                    0.0277093, 0.0409486,
                    0.0409486, 0.0643054,
                    0.0643054, 0.0755462,
                    0.0755462, 0.221729,
                    0.221729, 0.345984,
                    0.345984, 0.707055,
                    0.707055, 1.01989,
                    1.01989, 1.33125,
                    1.33125, 1.64993,
                    1.64993, 1.88383,
                    1.88383, 2.25367,
                    2.25367, 2.62643,
                    2.62643, 3.18193,
                    3.18193, 3.7842,
                    3.7842, 4.44202,
                    4.44202, 5.08084,
                    5.08084, 5.85414;



    } // End group size_cal


group: flow_cal {
    // Group containing calibration of flow rates of the PCASP
    //
    :title = "Flow calibration of PCASP";
    :comment = "Group containing sample flow calibration information. Sample flow output and/or input is measured by a calibrated meter";
    :references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp";

    // Define any group dimensions in addition to the global dimension, time.
    dimensions:
        max_flows = 1024;    // Maximum number of different flows in a calibration

    // Define group variables
    variables:
        string applies_to(time);
            applies_to:long_name = "Each calibration applies to these measurements";
            applies_to:comments = "String of applicable flight numbers for each calibration date";

        string traceability(time);
            traceability:long_name = "Traceability trail for each calibration";
            traceability:comment = "Link to file/s showing traceability of calibration materials and instruments";

        int cal_flag(time);
            cal_flag:long_name = "Flag denoting quality of calibration";
            cal_flag:valid_range = 0, 3;
            cal_flag:flag_values = 0, 1, 2, 3;
            cal_flag:flag_meanings = "good questionable poor missing_or_bad";
            cal_flag:_FillValue = 3;

        float flows_reported(time,max_flows);
            flows_reported:long_name = "Array of flow rates reported by PCASP for each value in flows_actual";
            flows_reported:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_reported for each time is the same as flows_actual for that time.";
            flows_reported:units = "cc/s";
            flows_reported:valid_min = 0;
            flows_reported:_FillValue = NaN;

        float flows_actual(time,max_flows);
            flows_actual:long_name = "Array of measured flow rate for each value in flows_reported";
            flows_actual:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_actual for each time is the same as flows_reported for that time.";
            flows_actual:units = "cc/s";
            flows_actual:valid_min = 0;
            flows_actual:_FillValue = NaN;

        string flow_fit(time);
            flow_fit:long_name = "Calibration equation of sample flow.";
            flow_fit:comment = "String of equation used to convert reported flow to calibrated flow rate. This will involve a fit to the data given for the same time stamp in the flows variable. A string is used for flexibility but may be changed to polynomial values in the future if appropriate.";
        flow_fit:_FillValue = "";
    

    data:
        // Data is comma-delineated with no additional deliniation between 
        // dimensions. Thus the data is presented flattened with the overall 
        // length being d1*d2*..dn. As specified in the variable definition,
        // the dimensions are cycled over in reverse order so for multi-
        // dimensional arrays, the last dimension varies fastest. Thus, 
        // row-order rather than column order is used for matrices.. If 
        // var = np.array([[11,12,13],[21,22,23]]) then var.flatten() or 
        // np.ravel(var) will write the array in the correct way.
    } // End group flow_cal

       

} // EOF