netcdf PCASP_faam_20191107_v001_r000_cal {

// global attributes:
		:Conventions = "CF-1.6" ;
		:institution = "FAAM. Facility for Airborne Atmospheric Measurements" ;
		:address = "Building 146, Cranfield University, Cranfield MK43 0AL UK" ;
		:title = "FAAM calibration data for the PCASP-2" ;
		:source = "Laboratory-based calibration" ;
		:instr = "PCASP-2" ;
		:instr_long_name = "Passive Cavity Spectrometer Probe. SPP200 electronics package" ;
		:instr_serialnumber = "PMI-1022-1202-31" ;
		:references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
		:username = "Graeme Nott <graeme.nott@faam.ac.uk>" ;
		:history = "20191202T1719 Initial creation" ;
		:software_version = "0.3" ;

group: bin_cal {
  dimensions:
  	time = UNLIMITED ; // (2 currently)
  	bin = 30 ;
  	bin_bounds = 2 ;
  variables:
  	float time(time) ;
  		time:standard_name = "time" ;
  		time:long_name = "time of calibration" ;
  		time:timezone = "UTC" ;
  		time:units = "days since 1970-01-01 00:00:00" ;
  		time:strftime_format = "days since %Y-%m-%d %Z" ;
  	int bin(bin) ;
  		bin:long_name = "bin number" ;
  		bin:comment = "The PCASP has 30 bins however the first has a somewhat undefined lower boundary and should therefore be discarded." ;
  	string applies_to(time) ;
  		applies_to:long_name = "Each calibration applies to these measurements" ;
  		applies_to:comment = "String of applicable flight numbers for calibration" ;
  	string descr(time) ;
  		descr:long_name = "Description of calibration" ;
  		descr:comment = "Campaign name/s for which these calibrations apply" ;
  	string traceability(time) ;
  		traceability:long_name = "Traceability trail for each calibration" ;
  		traceability:comment = "Unique lot numbers for each calibration PSL. These can be traced to the original NIST-traceable certificates." ;
  	int cal_flag(time) ;
  		cal_flag:long_name = "Flag denoting quality of calibration" ;
  		cal_flag:valid_range = 0, 3 ;
  		cal_flag:flag_values = 0, 1, 2, 3 ;
  		cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
  		cal_flag:_FillValue = 3 ;
  	int ADC_thres(time, bin, bin_bounds) ;
  		ADC_thres:long_name = "Lower and upper ADC thresholds for each bin" ;
  		ADC_thres:comment = "Coverage of each bin in terms of the digitized peak photovoltage. This variable has been included primarily for error checking as the same values should be in the standard data files." ;
  		ADC_thres:valid_range = 0, 1288 ;
  		ADC_thres:_FillValue = -2147483648 ;
  	float x-section(time, bin, bin_bounds) ;
  		x-section:long_name = "Scattering cross-section boundaries for each bin" ;
  		x-section:comment = "Lower boundary of first bin is undefined." ;
  		x-section:units = "m**2" ;
  		x-section:ancillary_variables = "x-section_width_err" ;
  		x-section:_FillValue = -9999.f ;
  	float x-section_err(time, bin, bin_bounds) ;
  		x-section_err:long_name = "Uncertainty of scattering cross section boundaries for each bin" ;
  		x-section_err:comment = "Straight-line fits for scattering cross-section versus ADC voltage are calculated along with sensitivities to the uncertainty in these data. See section 2.2.3 of Rosenberg et al. (2012) for details." ;
  		x-section_err:_FillValue = -9999.f ;
  	float x-section_width(time, bin) ;
  		x-section_width:long_name = "Width of each bin in terms of scattering cross section" ;
  	float x-section_width_err(time, bin) ;
  		x-section_width_err:long_name = "Uncertainty of scattering cross section boundaries for each bin" ;
  		x-section_width_err:comment = "" ;
  		x-section_width_err:flag_values = 0, 1 ;
  		x-section_width_err:flag_meanings = "Independent_uncertainties \n                                                 Dependent_uncertainties" ;
  		x-section_width_err:_FillValue = -9999.f ;
  	float dia_centre(time, bin) ;
  		dia_centre:long_name = "Centre diameter associated with each bin number for given particle material properties" ;
  		dia_centre:comment = "This is the weighted average of each of the regions of the scattering curve which include the range of scattering cross-sections in each bin with the uncertainty of these boundaries included. This is discussed in sections 4.1 and 4.2 of Rosenberg et al. (2012)." ;
  		dia_centre:refractive_index = "1.59+0i" ;
  		dia_centre:shape = "spherical" ;
  		dia_centre:units = "um" ;
  		dia_centre:ancillary_variables = "dia_centre_err dia_width" ;
  		dia_centre:_FillValue = -9999.f ;
  	float dia_centre_err(time, bin) ;
  		dia_centre_err:long_name = "Uncertainty of bin centre diameter" ;
  		dia_centre_err:comment = "See sections 4.1 and 4.2 of Rosenberg et al. (2012). for details." ;
  		dia_centre_err:units = "um" ;
  		dia_centre_err:_FillValue = -9999.f ;
  	float dia_width(time, bin) ;
  		dia_width:long_name = "Diameter width associated with each bin number for given particle material properties" ;
  		dia_width:comment = "This is the sum of all regions of the scattering curve which include the range of scattering cross-sections in each bin with the uncertainty of these boundaries included. This is discussed in sections 4.1 and 4.2 of Rosenberg et al. (2012)." ;
  		dia_width:refractive_index = "1.59+0i" ;
  		dia_width:shape = "spherical" ;
  		dia_width:units = "um" ;
  		dia_width:ancillary_variables = "dia_width_err" ;
  		dia_width:_FillValue = -9999.f ;
  	float dia_width_err(time, bin) ;
  		dia_width_err:long_name = "Uncertainty of bin width" ;
  		dia_width_err:comment = "See sections 4.1 and 4.2 of Rosenberg et al. (2012). for details." ;
  		dia_width_err:units = "um" ;
  		dia_width_err:_FillValue = -9999.f ;

  // group attributes:
  		:title = "Size bin calibration of PCASP" ;
  		:comment = "Group containing calibration of size bins of the PCASP. Photodetector voltage pulse-heights are calibrated to the calculated scattering cross-section of known PSL and DEHS monodisperse distributions. Data contained in this group is copied straight from the existing csv calibration files." ;
  		:references = "P.D. Rosenberg, A.R. Dean, P.I. Williams, J.R. Dorsey, A. Minikin, M.A. Pickering and A. Petzold, Particle sizing calibration with refractive index correction for light scattering optical particle counters and impacts upon PCASP and CDP data collected during the Fennec campaign, Atmos. Meas. Tech., 5, 1147-1163, doi:10.5194/amt-5-1147-2012, 2012." ;
  data:

   time = 18082, 18208 ;

   bin = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
      20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30 ;

   applies_to = _, _ ;

   descr = "ACRUISE-1. MOYA Arctic wetlands. ACSIS-5. ARNA-1", 
      "ACRUISE-1. MOYA Arctic wetlands. ACSIS-5. ARNA-1" ;

   traceability = 
      "125nm (#44245). 150nm (#202026). 203nm (#44793). 216nm (#16779). 240nm (#45059). 269nm (#166237). 303nm (#196947). 345nm (#199283). 400nm (#164245). 453nm (#166631). 508nm (#44115). 600nm (#166837). 707nm (#44582). 799nm (#164766). 903nm (#44869). 0.994um (#200992). 1.101um (#43973). 1.361um (#199629). 1.592um (#204268). 1.745um (#205235). 2.020um (#181058). 2.504um (#190272). 3.007um (#185943).", 
      "269nm (#166237). 303nm (#196947). 345nm (#199283). 400nm (#164245). 453nm (#166631). 508nm (#44115). 600nm (#166837). 707nm (#44582). 799nm (#164766). 903nm (#44869). 0.994um (#200992). 1.101um (#43973). 1.361um (#199629). 1.592um (#204268). 1.745um (#205235). 2.020um (#181058). 2.504um (#190272). 3.007um (#185943)." ;

   cal_flag = 1, 1 ;

   ADC_thres =
  20, 692,
  692, 1146,
  1146, 1814,
  1814, 2769,
  2769, 4096,
  4096, 4192,
  4192, 4231,
  4231, 4282,
  4282, 4348,
  4348, 4537,
  4537, 4825,
  4825, 5251,
  5251, 5859,
  5859, 6703,
  6703, 8192,
  8192, 8335,
  8335, 8435,
  8435, 8520,
  8520, 8767,
  8767, 8981,
  8981, 9194,
  9194, 9412,
  9412, 9572,
  9572, 9825,
  9825, 10080,
  10080, 10460,
  10460, 10872,
  10872, 11322,
  11322, 11759,
  11759, 12288,
  20, 692,
  692, 1146,
  1146, 1814,
  1814, 2769,
  2769, 4096,
  4096, 4192,
  4192, 4231,
  4231, 4282,
  4282, 4348,
  4348, 4537,
  4537, 4825,
  4825, 5251,
  5251, 5859,
  5859, 6703,
  6703, 8192,
  8192, 8335,
  8335, 8435,
  8435, 8520,
  8520, 8767,
  8767, 8981,
  8981, 9194,
  9194, 9412,
  9412, 9572,
  9572, 9825,
  9825, 10080,
  10080, 10460,
  10460, 10872,
  10872, 11322,
  11322, 11759,
  11759, 12288 ;

   x-section =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

   x-section_err =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

   x-section_width =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _ ;

   x-section_width_err =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _ ;

   dia_centre =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _ ;

   dia_centre_err =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _ ;

   dia_width =
  _, _, _, _, _, _, 0.00119786, 0.00156644, 0.00202715, 0.00580503, 
      0.00884576, 0.0130844, 0.0186744, 0.025923, 0.0457338, 0.359616, 
      0.255995, 0.217595, 0.632307, 0.547828, 0.545268, 0.558068, 0.409591, 
      0.647666, 0.652786, 0.972779, 1.0547, 1.15198, 1.1187, 1.35421,
  _, _, _, _, _, _, 0.000882833, 0.00115447, 0.00149403, 0.00427835, 
      0.00651938, 0.00964326, 0.0137631, 0.0191054, 0.0337061, 0.266736, 
      0.185376, 0.15757, 0.457879, 0.396705, 0.394852, 0.40412, 0.296602, 
      0.469002, 0.47271, 0.70443, 0.76375, 0.834193, 0.810094, 0.980641 ;

   dia_width_err =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _ ;
  } // group bin_cal

group: flow_cal {
  dimensions:
  	time = UNLIMITED ; // (1 currently)
  	max_flows = 1024 ;
  variables:
  	float time(time) ;
  		time:standard_name = "time" ;
  		time:long_name = "time of calibration" ;
  		time:timezone = "UTC" ;
  		time:units = "days since 1970-01-01 00:00:00" ;
  		time:strftime_format = "days since %Y-%m-%d %Z" ;
  	string applies_to(time) ;
  		applies_to:long_name = "Each calibration applies to these measurements" ;
  		applies_to:comments = "String of applicable flight numbers for calibration" ;
  	string descr(time) ;
  		descr:long_name = "Description of calibration" ;
  		descr:comment = "Campaign name/s for which these calibrations apply" ;
  	string traceability(time) ;
  		traceability:long_name = "Traceability trail for each calibration" ;
  		traceability:comment = "Calibration of low flow cell s/n 1702010-L" ;
  	int cal_flag(time) ;
  		cal_flag:long_name = "Flag denoting quality of calibration" ;
  		cal_flag:valid_range = 0, 3 ;
  		cal_flag:flag_values = 0, 1, 2, 3 ;
  		cal_flag:flag_meanings = "good questionable poor missing_or_bad" ;
  		cal_flag:_FillValue = 3 ;
  	float flows_reported(time, max_flows) ;
  		flows_reported:long_name = "Array of flow rates reported by PCASP for each value in flows_actual" ;
  		flows_reported:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_reported for each time is the same as flows_actual for that time." ;
  		flows_reported:units = "cc/s" ;
  		flows_reported:_FillValue = NaNf ;
  	float flows_actual(time, max_flows) ;
  		flows_actual:long_name = "Array of actual flow rates for each value in flows_reported" ;
  		flows_actual:comment = "The number of different flows included in each calibration will differ depending on operator and circumstance. The maximum possible flows is given by the dimension max_flows. The variable is padded by the _FillValue. It is the users obligation to check that the number of flows_actual for each time is the same as flows_reported for that time." ;
  		flows_actual:units = "cc/s" ;
  		flows_actual:_FillValue = NaNf ;
  	string flow_fit(time) ;
  		flow_fit:long_name = "Calibration equation of sample flow." ;
  		flow_fit:comment = "String of equation used to convert reported flow to calibrated flow rate. This will involve a fit to the data given for the same time stamp in the flows variable. A string is used for flexibility but may be changed to polynomial values in the future if appropriate." ;
  		string flow_fit:_FillValue = "" ;

  // group attributes:
  		:title = "Flow calibration of PCASP" ;
  		:comment = "Gilibrator 2 small cell (to 250cc/m) connected to outlet of PCASP1. Small CV needle valve used to throttle inlet flow with inline Alicat flowmeter used to measure T & P of inlet air" ;
  		:references = "http://www.faam.ac.uk/index.php/science-instruments/aerosol/304-pcasp" ;
  data:

   time = 17660 ;

   applies_to = "C173-" ;

   descr = _ ;

   traceability = 
      "Calibrated 20170210. Uncertainty of flow = 0.44% + instrument resolution." ;

   cal_flag = 0 ;

   flows_reported =
  1.046, 0.996, 0.911, 0.789, 0.72, 0.611, 0.522, 0.397, 0.334, 0.235, 
      0.148, 0.115, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _ ;

   flows_actual =
  0.919, 0.879, 0.808, 0.699, 0.64, 0.542, 0.455, 0.344, 0.275, 0.185, 
      0.071, 0.022, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _, _, _, _, _, _ ;

   flow_fit = "0.280*x**3 - 0.672*x**2 + 1.397*x - 0.123" ;
  } // group flow_cal
}
